
package mem_pkg;

  import uvm_pkg::*;

  `include "mem.svh"
  `include "mem_seq_lib.svh"

endpackage : mem_pkg

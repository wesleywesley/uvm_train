
package test_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import packet_pkg::*;
  import datain_agt_pkg::*;

  `include "agent_test.svh"

  `include "anlsp.svh"
  `include "anlsp_test.svh"

  `include "my_hello_world.svh"
  `include "triple.svh"

endpackage : test_pkg

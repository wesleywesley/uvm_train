
package switch_model_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import mem_pkg::*;
  import packet_pkg::*;
  import datain_agt_pkg::*;
  import dataout_agt_pkg::*;
  import mem_agt_pkg::*;
  
  `include "switch_model.svh"

endpackage : switch_model_pkg

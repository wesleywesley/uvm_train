
package switch_env_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import mem_pkg::*;
  import packet_pkg::*;
  import datain_agt_pkg::*;
  import dataout_agt_pkg::*;
  import mem_agt_pkg::*;
  import switch_env_pkg::*;
  
  `include "switch_env.svh"

endpackage : switch_env_pkg

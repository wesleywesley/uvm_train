
package packet_pkg;

  import uvm_pkg::*;

  `include "packet.svh"
  `include "packet_seq_lib.svh"

endpackage : packet_pkg
